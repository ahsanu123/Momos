CircuitMaker Text
5.6
Probes: 3
U1_6
Transient Analysis
0 633 143 65280
V4_1
Transient Analysis
1 465 153 65535
U1_6
AC Analysis
0 626 146 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
40 0 30 150 10
176 80 1364 747
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
27 D:\CircuitMaker2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 1532 509
9961490 0
0
6 Title:
5 Name:
0
0
0
11
2 +V
167 531 222 0 1 3
0 3
0
0 0 54256 180
2 1v
7 -2 21 6
2 V1
7 -12 21 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3409 0 0
2
44951 0
0
7 Ground~
168 465 107 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3951 0 0
2
44951 0
0
7 Ground~
168 466 177 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8885 0 0
2
44951 0
0
11 Signal Gen~
195 419 157 0 19 64
0 6 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1186693120 0 1065353216
20
1 24000 0 1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
5 -1/1V
-18 -30 17 -22
2 V4
-7 -40 7 -32
0
0
37 %D %1 %2 DC 0 SIN(0 1 24k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
3780 0 0
2
44951 0
0
10 Op-Amp5:A~
219 568 145 0 5 11
0 7 5 8 2 4
0
0 0 848 692
8 LM358/NS
16 -25 72 -17
2 U1
37 -35 51 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
0
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 0 0 0 0 0
1 U
9265 0 0
2
44951 3
0
2 +V
167 568 187 0 1 3
0 8
0
0 0 53616 180
2 5V
7 -7 21 1
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
9442 0 0
2
44951 2
0
7 Ground~
168 568 119 0 1 3
0 2
0
0 0 53360 180
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9424 0 0
2
44951 1
0
9 Resistor~
219 593 91 0 2 5
0 5 4
0
0 0 880 0
4 2.2k
-14 -14 14 -6
2 R6
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 48249868
82 0 0 0 1 0 0 0
1 R
9968 0 0
2
44951 0
0
9 Resistor~
219 510 91 0 3 5
0 2 5 -1
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R5
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 250
82 0 0 0 1 0 0 0
1 R
9281 0 0
2
44951 0
0
9 Resistor~
219 493 152 0 2 5
0 6 7
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 38741340
82 0 0 0 1 0 0 0
1 R
8464 0 0
2
44951 0
0
9 Resistor~
219 531 187 0 3 5
0 3 7 1
0
0 0 880 90
2 1k
9 0 23 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7168 0 0
2
44951 0
0
11
1 1 3 0 0 4224 0 1 11 0 0 2
531 207
531 205
5 2 4 0 0 4224 0 5 8 0 0 4
586 145
653 145
653 91
611 91
1 1 2 0 0 8320 0 2 9 0 0 3
465 101
465 91
492 91
2 0 5 0 0 8320 0 5 0 0 5 3
550 139
541 139
541 91
1 2 5 0 0 0 0 8 9 0 0 2
575 91
528 91
1 2 2 0 0 16 0 3 4 0 0 3
466 171
466 162
450 162
1 1 6 0 0 4224 0 4 10 0 0 2
450 152
475 152
2 0 7 0 0 4224 0 10 0 0 9 2
511 152
531 152
2 1 7 0 0 0 0 11 5 0 0 3
531 169
531 151
550 151
1 4 2 0 0 0 0 7 5 0 0 2
568 127
568 132
1 3 8 0 0 4224 0 6 5 0 0 2
568 172
568 158
0
0
8 0 0
0
0
0
0 0 0
0
0 0 0
1000 1 1 500000
0 0.0002083 8.333e-07 8.333e-07
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
