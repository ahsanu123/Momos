CircuitMaker Text
5.6
Probes: 3
U1_6
AC Analysis
0 639 181 65280
V2_1
AC Analysis
1 154 176 65535
U2_6
Transient Analysis
0 338 172 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 405
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
27 D:\CircuitMaker2000\BOM.DAT
0 7
2 2 0.500000 0.500000
344 176 1532 509
9961490 0
0
6 Title:
5 Name:
0
0
0
19
7 Ground~
168 628 307 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5130 0 0
2
44951.2 0
0
10 Capacitor~
219 516 211 0 2 5
0 2 7
0
0 0 848 90
5 470pF
-50 -5 -15 3
2 C1
-28 -14 -14 -6
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
391 0 0
2
44951.2 0
0
10 Capacitor~
219 527 117 0 2 5
0 9 4
0
0 0 848 0
7 0.001uF
-24 -18 25 -10
2 C2
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3124 0 0
2
44951.2 1
0
7 Ground~
168 516 235 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3421 0 0
2
44951.2 2
0
7 Ground~
168 591 216 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8157 0 0
2
44951.2 3
0
2 +V
167 591 146 0 1 3
0 8
0
0 0 53616 0
2 15
-7 -22 7 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5572 0 0
2
44951.2 4
0
10 Op-Amp5:A~
219 591 181 0 5 11
0 7 3 8 2 4
0
0 0 848 0
8 LM358/NS
16 -25 72 -17
2 U1
37 -35 51 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
0
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 0 1 0 0 0
1 U
8901 0 0
2
44951.2 5
0
2 +V
167 262 219 0 1 3
0 10
0
0 0 53616 180
2 5V
7 -7 21 1
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7361 0 0
2
5.90063e-315 0
0
7 Ground~
168 262 139 0 1 3
0 2
0
0 0 53360 180
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4747 0 0
2
5.90063e-315 5.26354e-315
0
2 +V
167 214 266 0 1 3
0 12
0
0 0 54256 180
2 1v
7 -2 21 6
2 V3
7 -12 21 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
972 0 0
2
5.90063e-315 5.30499e-315
0
10 Op-Amp5:A~
219 262 173 0 5 11
0 6 5 10 2 5
0
0 0 848 692
8 LM358/NS
16 -25 72 -17
2 U2
37 -35 51 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
0
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 0 1 0 0 0
1 U
3472 0 0
2
5.90063e-315 5.32571e-315
0
7 Ground~
168 146 204 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9998 0 0
2
5.90063e-315 5.34643e-315
0
11 Signal Gen~
195 101 184 0 64 64
0 11 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1176256512 0 1065353216
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
1 10000 0 1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
5 -1/1V
-18 -30 17 -22
2 V2
-7 -40 7 -32
0
0
37 %D %1 %2 DC 0 SIN(0 1 10k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3536 0 0
2
5.90063e-315 5.3568e-315
0
9 Resistor~
219 628 269 0 3 5
0 2 3 -1
0
0 0 880 90
3 10k
5 0 26 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 22
82 0 0 0 1 0 0 0
1 R
4597 0 0
2
44951.2 0
0
9 Resistor~
219 628 218 0 2 5
0 3 4
0
0 0 880 90
3 22k
5 0 26 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 80882360
82 0 0 0 1 0 0 0
1 R
3835 0 0
2
44951.2 0
0
9 Resistor~
219 413 175 0 2 5
0 5 9
0
0 0 880 0
4 9.1k
-13 -14 15 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3670 0 0
2
44951.2 6
0
9 Resistor~
219 492 175 0 2 5
0 9 7
0
0 0 880 0
4 6.2k
-14 -14 14 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5616 0 0
2
44951.2 7
0
9 Resistor~
219 177 179 0 2 5
0 11 6
0
0 0 880 0
3 100
-10 -14 11 -6
2 R6
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 62
82 0 0 0 1 0 0 0
1 R
9323 0 0
2
5.90063e-315 5.36716e-315
0
9 Resistor~
219 214 218 0 3 5
0 12 6 1
0
0 0 880 90
3 100
5 0 26 8
2 R5
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 250
82 0 0 0 1 0 0 0
1 R
317 0 0
2
5.90063e-315 5.37752e-315
0
21
0 2 3 0 0 4224 0 0 7 3 0 4
628 247
565 247
565 187
573 187
1 1 2 0 0 4096 0 1 14 0 0 2
628 301
628 287
2 1 3 0 0 0 0 14 15 0 0 2
628 251
628 236
2 0 4 0 0 4096 0 15 0 0 9 2
628 200
628 181
1 0 5 0 0 8192 0 16 0 0 8 4
395 175
395 174
336 174
336 173
2 0 6 0 0 4096 0 19 0 0 7 2
214 200
214 179
2 1 6 0 0 4224 0 18 11 0 0 2
195 179
244 179
2 5 5 0 0 12416 0 11 11 0 0 6
244 167
236 167
236 116
336 116
336 173
280 173
2 5 4 0 0 4224 0 3 7 0 0 4
536 117
673 117
673 181
609 181
2 0 7 0 0 4096 0 2 0 0 11 2
516 202
516 175
1 2 7 0 0 4224 0 7 17 0 0 2
573 175
510 175
1 4 2 0 0 4224 0 5 7 0 0 2
591 210
591 194
1 3 8 0 0 4224 0 6 7 0 0 2
591 155
591 168
1 1 2 0 0 0 0 4 2 0 0 2
516 229
516 220
1 0 9 0 0 4224 0 3 0 0 16 3
518 117
453 117
453 175
1 2 9 0 0 0 0 17 16 0 0 2
474 175
431 175
1 3 10 0 0 4224 0 8 11 0 0 4
262 204
262 184
262 184
262 186
1 4 2 0 0 0 0 9 11 0 0 2
262 147
262 160
1 1 11 0 0 4224 0 18 13 0 0 2
159 179
132 179
1 1 12 0 0 4224 0 10 19 0 0 2
214 251
214 236
1 2 2 0 0 0 0 12 13 0 0 3
146 198
146 189
132 189
0
0
17 0 0
0
0
0
0 0 0
0
0 0 0
600 1 1 40000
0 0.001 8.333e-07 8.333e-07
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
